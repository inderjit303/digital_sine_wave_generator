* /home/inderjitsingh/eSim_Mixed_signal_marathon_2022/counter_4b/counter_4b.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat 05 Mar 2022 12:50:47 PM UTC

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ inderjit_4bitcounter		
U11  ? ? ? ? adc_bridge_2		
U5  clk reset Net-_U2-Pad1_ Net-_U2-Pad2_ adc_bridge_2		
U6  Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_R3-Pad1_ o2 o1 o0 dac_bridge_4		
R3  Net-_R3-Pad1_ o3 1k		
C1  o3 GND 1u		
v1  Net-_R1-Pad1_ GND pulse		
v3  ? ? pulse		
v2  reset GND pulse		
R1  Net-_R1-Pad1_ clk 1k		
R2  clk GND 1k		
U1  ? plot_v1		
U10  o3 plot_v1		
U7  o2 plot_v1		
U8  o1 plot_v1		
U9  o0 plot_v1		
U3  reset plot_v1		
U4  clk plot_v1		

.end
