* /home/inderjitsingh/eSim_Mixed_signal_marathon_2022/digital_sine_wave/digital_sine_wave.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu 10 Mar 2022 09:46:53 AM UTC

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ inderjit_prs8bit_generator		
U2  Net-_U2-Pad1_ Net-_U1-Pad3_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U2-Pad7_ Net-_U2-Pad8_ Net-_U2-Pad9_ Net-_U2-Pad10_ inderjit_digi_sinewave_generator		
U3  clk reset Net-_U1-Pad1_ Net-_U1-Pad2_ adc_bridge_2		
U6  Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U2-Pad7_ Net-_U2-Pad8_ Net-_U2-Pad9_ Net-_U2-Pad10_ Net-_U6-Pad9_ Net-_U6-Pad10_ Net-_U6-Pad11_ Net-_U6-Pad12_ Net-_U6-Pad13_ Net-_U6-Pad14_ Net-_U6-Pad15_ Net-_U6-Pad16_ dac_bridge_8		
v1  clk GND pulse		
v2  reset GND pulse		
R1  dac_out Net-_L1-Pad1_ 130		
U7  dac_out plot_v1		
U8  analog_out plot_v1		
U4  reset plot_v1		
U5  clk plot_v1		
L1  Net-_L1-Pad1_ analog_out 10mH		
C2  analog_out GND 2.5u		
X1  Net-_U6-Pad16_ Net-_U6-Pad15_ Net-_U6-Pad14_ Net-_U6-Pad13_ Net-_U6-Pad12_ Net-_U6-Pad11_ Net-_U6-Pad10_ Net-_U6-Pad9_ GND GND dac_out 10bitDAC		
U9  clk Net-_U2-Pad1_ adc_bridge_1		

.end
